//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// System-Verilog Alex Grinshpun May 2018
// New coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering 2019 


module	step_controller	(
					input		logic	clk,
					input		logic	resetN,
					input 	logic	[10:0] pixelX,// current VGA pixel 
					input 	logic	[10:0] pixelY,
					
					output	logic [2:0] step_type,
					output 	logic	[10:0] tileTopLeftX, 
					output 	logic	[10:0] tileTopLeftY,
					output	logic	drawingRequest, // indicates pixel inside the bracket
					output	logic	[7:0]	 RGBout //optional color output for mux 
);

//__________________________________
parameter  int Tile_WIDTH_X = 6; // 2^6=64
parameter  int Tile_HEIGHT_Y = 6;// 2^6=64
//__________________________________
const logic [2:0] FREE=3'b000, REGULAR_STEP=3'b001;
//parameter  int NUM_OF_ROWS = 7;
//parameter  int NUM_OF_COLS = 10;

parameter  logic [7:0] OBJECT_COLOR = 8'h5b; 

/*
logic [0:2] [0:2] [2:0] tile_map = {
{REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP},
{FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE},
{FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE},
{FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE},
{FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE},
{FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE},
{FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE}, //Not Used
{FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE}  //Not Used
};
*/

parameter  int BRICK_WIDTH_X = 16;
parameter  int BRICK_HEIGHT_Y = 16;

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// bitmap  representation for a transparent pixel 

parameter  int NUM_OF_ROWS = 30;
parameter  int NUM_OF_COLS = 30;

const logic [0:NUM_OF_COLS-1] [0:NUM_OF_ROWS-1] [1:0] tile_map = {
	{REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP},
	{REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,FREE,FREE,FREE,FREE,FREE,FREE,REGULAR_STEP,REGULAR_STEP,FREE,FREE,FREE,REGULAR_STEP},
	{REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP,REGULAR_STEP}
};

// Frame size
const int x_FRAME_SIZE = 639 ;
const int y_FRAME_SIZE = 479 ;

const int x_GRID_SIZE = y_FRAME_SIZE;
const int y_GRID_SIZE = y_FRAME_SIZE;

int X_index_in_grid ; 
int X_index_in_grid_delayed ; 
int y_index_in_grid ;
logic	[10:0] topLeftY;
logic inside_grid;
//logic	[10:0] X_VGA_DELAY = x_vga_delay_debug;
const logic [10:0] x_vga_delay_debug = 2;
assign X_index_in_grid = ((pixelX)>> 4);
assign X_index_in_grid_delayed = ((pixelX - x_vga_delay_debug )>> 4);
assign y_index_in_grid = (pixelY >> 4);
assign inside_grid = (pixelX <= x_GRID_SIZE);

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN)
	begin
		RGBout			<=	8'b0;
		drawingRequest	<=	0;
	end
	else
	begin
		
		//drawing offset logic
		if (inside_grid ) // test if it is inside the grid (int a delay of some clocks)
		begin 
			RGBout  <= OBJECT_COLOR ;	// colors table 
			//draw logic
			drawingRequest <= (tile_map[y_index_in_grid][X_index_in_grid] == REGULAR_STEP) ;
			tileTopLeftX	<= (pixelX % BRICK_WIDTH_X); //calculate relative offsets from top left corner of the brick
			tileTopLeftY	<= (pixelY % BRICK_HEIGHT_Y); //calculate relative offsets from top left corner of the brick
		end 
		else
		begin  
			RGBout <= TRANSPARENT_ENCODING ; // so it will not be displayed 
			drawingRequest <= 1'b0 ;// transparent color 
			tileTopLeftX	<= 0; //no offset
			tileTopLeftY	<= 0; //no offset
		end 
	end
end 





/*
assign step_type = tile_map[pixelY >> Tile_HEIGHT_Y][pixelX >> Tile_WIDTH_X];
assign tileTopLeftX = (pixelX >> Tile_WIDTH_X) << Tile_WIDTH_X;
assign tileTopLeftY = (pixelY >> Tile_HEIGHT_Y) << Tile_HEIGHT_Y;



always_ff@(posedge clk)
begin
	if(tile_map[pixelY >> Tile_HEIGHT_Y][pixelX >> Tile_WIDTH_X] == REGULAR_STEP) begin
		RGBout  <= OBJECT_COLOR;
		drawingRequest <= 1'b1;
	end
	step_type <= tile_map[pixelY >> Tile_HEIGHT_Y][pixelX >> Tile_WIDTH_X];
	tileTopLeftX <= (pixelX >> Tile_WIDTH_X) << Tile_WIDTH_X;
	tileTopLeftY <= (pixelY >> Tile_HEIGHT_Y) << Tile_HEIGHT_Y;
end 

*/

endmodule
