
module	buttons_bitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input	logic [2:0] button_type,
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 7;  // 2^7 = 128
localparam  int OBJECT_NUMBER_OF_X_BITS = 7;  // 2^7 = 128 


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;

// generating a smiley bitmap

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h2F ;// RGB value in the bitmap representing a transparent pixel 

logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {
{8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h00, 8'h00, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hFA, 8'hFA, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hFA, 8'hFA, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hFA, 8'hFA, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h88, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'hFA, 8'hFA, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h24, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h20, 8'h64, 8'h64, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h24, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h20, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h00, 8'h00, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h44, 8'h88, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hFA, 8'hFA, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h64, 8'h64, 8'h64, 8'h64, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h49, 8'h49, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h49, 8'h49, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h49, 8'h49, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hDB, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'hDB, 8'hDB, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'hDB, 8'hDB, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'hDB, 8'hDB, 8'h92, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h04, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h04, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h04, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h04, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h04, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h04, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h92, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h00, 8'h00, 8'h04, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h6D, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h49, 8'h49, 8'h49, 8'h49, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h49, 8'h49, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F },
{8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F, 8'h2F }
};

// pipeline (ff) to get the pixel color from the array 	 

//////////--------------------------------------------------------------------------------------------------------------=

const logic [2:0] FREE=3'b000, REGU=3'b001, SLCT=3'b010;

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		if (InsideRectangle == 1'b1 )  // inside an external bracket 
			case(button_type)
				REGU: begin
					RGBout <= object_colors[offsetY+50][offsetX];
				end
				SLCT:begin
					RGBout <= object_colors[offsetY][offsetX];
				end
			endcase
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule