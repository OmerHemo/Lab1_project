
module	regular_step_bitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input	logic [2:0] step_type,
					input	logic [2:0] brake_state,
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 6;  // 2^6 = 64 
localparam  int OBJECT_NUMBER_OF_X_BITS = 6;  // 2^4 = 64 


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;

// generating a smiley bitmap

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h13 ;// RGB value in the bitmap representing a transparent pixel 

logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'hB0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'h13, 8'hE0, 8'hE0, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'hE0, 8'h13, 8'hE0, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'hE0, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hC8, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'h88, 8'hC8, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'h88, 8'hC8, 8'h88, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'h88, 8'hE0, 8'hE0, 8'hC8, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h88, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'h88, 8'hC8, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'h88, 8'hE0, 8'hE0, 8'hC8, 8'hE0, 8'hE0, 8'h88, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h00, 8'h88, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'h88, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'h88, 8'hE0, 8'h88, 8'hE0, 8'h88, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'h88, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'hE0, 8'h88, 8'hC8, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'h88, 8'hE0, 8'hC8, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h88, 8'h88, 8'hE0, 8'h88, 8'hE0, 8'h88, 8'h88, 8'h88, 8'hC8, 8'h88, 8'hE0, 8'hE0, 8'hE0, 8'h88, 8'h88, 8'hC8, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'hE0, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'hE0, 8'h13, 8'h13, 8'hE0, 8'hE0, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h97, 8'h97, 8'h49, 8'h97, 8'h97, 8'h97, 8'h49, 8'h49, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h49, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h49, 8'h49, 8'h49, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hE8, 8'h97, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'h97, 8'hE8, 8'h49, 8'hE8, 8'h49, 8'h49, 8'h97, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'h49, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'h49, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'h49, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h97, 8'h97, 8'h49, 8'h49, 8'h49, 8'h97, 8'h49, 8'h49, 8'h97, 8'h97, 8'h49, 8'h97, 8'h97, 8'h97, 8'h97, 8'h49, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h49, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h49, 8'h49, 8'h97, 8'h49, 8'h97, 8'h49, 8'h49, 8'h49, 8'h97, 8'h97, 8'h49, 8'h97, 8'h97, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'h49, 8'h49, 8'h49, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h49, 8'hE8, 8'h97, 8'h49, 8'hE8, 8'h49, 8'h49, 8'hE8, 8'h49, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'h49, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'h49, 8'h49, 8'hE8, 8'hE8, 8'hE8, 8'h97, 8'hE8, 8'hE8, 8'hE8, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h5C, 8'h5C, 8'h0C, 8'h0C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h0C, 8'h0C, 8'h5C, 8'h5C, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h5C, 8'h5C, 8'h0C, 8'h0C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h0C, 8'h0C, 8'h5C, 8'h5C, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'h5C, 8'h5C, 8'h0C, 8'h0C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h0C, 8'h0C, 8'h5C, 8'h5C, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h00, 8'h5C, 8'h0C, 8'h0C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h5C, 8'h0C, 8'h0C, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'h00, 8'hFF, 8'hDF, 8'hDF, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'h00, 8'h00, 8'h00, 8'h13, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hDF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDF, 8'hDF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDF, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hDF, 8'hDF, 8'hDF, 8'h00, 8'h00, 8'h13, 8'h00, 8'h00, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h00, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h00, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hFF, 8'hF0, 8'hF0, 8'hF0, 8'hFF, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hFF, 8'hFF, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h00, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h00, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hFF, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 },
{8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13 }
};

// pipeline (ff) to get the pixel color from the array 	 

//////////--------------------------------------------------------------------------------------------------------------=

const logic [2:0] FREE=3'b000, REGU=3'b001, GATE=3'b010, COIN=3'b011, PORT=3'b100, SPIK=3'b101, BRAK=3'b110;
const logic	[10:0] size_of_sep_y = 7;

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		if (InsideRectangle == 1'b1 )  // inside an external bracket 
			case(step_type)
				REGU: begin
					RGBout <= object_colors[offsetY][offsetX];
				end
				SPIK:begin
					RGBout <= object_colors[offsetY + 7][offsetX];
				end
				BRAK:begin
					case(brake_state)
						3:begin
							RGBout <= object_colors[offsetY + 14][offsetX];
						end
						2:begin
							RGBout <= object_colors[offsetY + 21][offsetX];
						end
						1:begin
							RGBout <= object_colors[offsetY + 28][offsetX];
						end
					endcase
				end
				PORT:begin
					RGBout <= object_colors[offsetY + 35][offsetX];
				end
				GATE:begin
					RGBout <= object_colors[offsetY + 42][offsetX];
				end
				COIN:begin
					RGBout <= object_colors[offsetY + 49][offsetX];
				end
			endcase
			//RGBout <= object_colors[offsetY][offsetX];	 
			//RGBout <=  {HitEdgeCode, 4'b0000 } ;  //get RGB from the colors table, option  for debug 
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule